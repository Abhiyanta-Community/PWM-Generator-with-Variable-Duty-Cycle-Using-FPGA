library verilog;
use verilog.vl_types.all;
entity pwm_5_variation_vlg_vec_tst is
end pwm_5_variation_vlg_vec_tst;
