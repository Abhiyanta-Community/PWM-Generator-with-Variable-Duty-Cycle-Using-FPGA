library verilog;
use verilog.vl_types.all;
entity pwm_5_variation_vlg_check_tst is
    port(
        \out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pwm_5_variation_vlg_check_tst;
